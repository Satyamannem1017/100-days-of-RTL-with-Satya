module add_sub(input [3:0]a,b,input m,output 
