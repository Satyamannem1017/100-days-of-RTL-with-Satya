`timescale 1ns/1ps
module clock(clk)
  input clk;
endmodule
